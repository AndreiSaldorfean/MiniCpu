-- Test bench script
library ieee;
use ieee.std_logic_1164.all; --include arrays

entity alu_tb is

end alu_tb;

architecture alu_arch_tb of alu_tb is

begin

end alu_arch_tb;