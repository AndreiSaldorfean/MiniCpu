library ieee;
use ieee.std_logic_1164.all; --include arrays

entity alu_entity is

end alu_entity;

architecture alu_arch of alu_entity is

begin

end alu_arch;